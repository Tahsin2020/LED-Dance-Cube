// UART_comp.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module UART_comp (
		input  wire  clk_clk,       //      clk.clk
		input  wire  gpio_035_rxd,  // gpio_035.rxd
		output wire  gpio_035_txd,  //         .txd
		input  wire  reset_reset_n  //    reset.reset_n
	);

	wire  [15:0] uart_custom_component_0_avm_m0_readdata;    // mm_interconnect_0:UART_custom_component_0_avm_m0_readdata -> UART_custom_component_0:avm_m0_readdata
	wire         uart_custom_component_0_avm_m0_waitrequest; // mm_interconnect_0:UART_custom_component_0_avm_m0_waitrequest -> UART_custom_component_0:avm_m0_waitrequest
	wire   [7:0] uart_custom_component_0_avm_m0_address;     // UART_custom_component_0:avm_m0_address -> mm_interconnect_0:UART_custom_component_0_avm_m0_address
	wire         uart_custom_component_0_avm_m0_read;        // UART_custom_component_0:avm_m0_read -> mm_interconnect_0:UART_custom_component_0_avm_m0_read
	wire         uart_custom_component_0_avm_m0_write;       // UART_custom_component_0:avm_m0_write -> mm_interconnect_0:UART_custom_component_0_avm_m0_write
	wire  [15:0] uart_custom_component_0_avm_m0_writedata;   // UART_custom_component_0:avm_m0_writedata -> mm_interconnect_0:UART_custom_component_0_avm_m0_writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;     // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;       // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;        // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;           // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;  // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;          // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;      // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         rst_controller_reset_out_reset;             // rst_controller:reset_out -> [UART_custom_component_0:reset_reset, mm_interconnect_0:UART_custom_component_0_reset_reset_bridge_in_reset_reset, uart_0:reset_n]

	new_component uart_custom_component_0 (
		.avm_m0_address     (uart_custom_component_0_avm_m0_address),     // avm_m0.address
		.avm_m0_read        (uart_custom_component_0_avm_m0_read),        //       .read
		.avm_m0_readdata    (uart_custom_component_0_avm_m0_readdata),    //       .readdata
		.avm_m0_write       (uart_custom_component_0_avm_m0_write),       //       .write
		.avm_m0_writedata   (uart_custom_component_0_avm_m0_writedata),   //       .writedata
		.avm_m0_waitrequest (uart_custom_component_0_avm_m0_waitrequest), //       .waitrequest
		.clock_clk          (clk_clk),                                    //  clock.clk
		.reset_reset        (rst_controller_reset_out_reset)              //  reset.reset
	);

	UART_comp_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (gpio_035_rxd),                              // external_connection.export
		.txd           (gpio_035_txd),                              //                    .export
		.irq           ()                                           //                 irq.irq
	);

	UART_comp_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                             (clk_clk),                                    //                                           clk_0_clk.clk
		.UART_custom_component_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),             // UART_custom_component_0_reset_reset_bridge_in_reset.reset
		.UART_custom_component_0_avm_m0_address                    (uart_custom_component_0_avm_m0_address),     //                      UART_custom_component_0_avm_m0.address
		.UART_custom_component_0_avm_m0_waitrequest                (uart_custom_component_0_avm_m0_waitrequest), //                                                    .waitrequest
		.UART_custom_component_0_avm_m0_read                       (uart_custom_component_0_avm_m0_read),        //                                                    .read
		.UART_custom_component_0_avm_m0_readdata                   (uart_custom_component_0_avm_m0_readdata),    //                                                    .readdata
		.UART_custom_component_0_avm_m0_write                      (uart_custom_component_0_avm_m0_write),       //                                                    .write
		.UART_custom_component_0_avm_m0_writedata                  (uart_custom_component_0_avm_m0_writedata),   //                                                    .writedata
		.uart_0_s1_address                                         (mm_interconnect_0_uart_0_s1_address),        //                                           uart_0_s1.address
		.uart_0_s1_write                                           (mm_interconnect_0_uart_0_s1_write),          //                                                    .write
		.uart_0_s1_read                                            (mm_interconnect_0_uart_0_s1_read),           //                                                    .read
		.uart_0_s1_readdata                                        (mm_interconnect_0_uart_0_s1_readdata),       //                                                    .readdata
		.uart_0_s1_writedata                                       (mm_interconnect_0_uart_0_s1_writedata),      //                                                    .writedata
		.uart_0_s1_begintransfer                                   (mm_interconnect_0_uart_0_s1_begintransfer),  //                                                    .begintransfer
		.uart_0_s1_chipselect                                      (mm_interconnect_0_uart_0_s1_chipselect)      //                                                    .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
