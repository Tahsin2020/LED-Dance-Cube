
module UART_comp (
	clk_clk,
	gpio_035_rxd,
	gpio_035_txd,
	reset_reset_n);	

	input		clk_clk;
	input		gpio_035_rxd;
	output		gpio_035_txd;
	input		reset_reset_n;
endmodule
